module Gaussian_Filter(


);
