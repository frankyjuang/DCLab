// (19 * 28) * 3 = 1596
parameter [32:0] COEF [1595:0] = '{
5442,367,5245,5342,451,5186,5205,460,5245,5167,281,5223,5064,325,5199,4945,355,5207,4833,376,5214,4782,176,5194,4669,181,5244,4578,197,5200,4491,180,5232,4377,234,5208,4290,243,5198,4161,252,5207,4117,250,5207,3988,239,5198,3901,221,5187,3770,221,5189,3704,209,5189,3590,174,5223,3499,165,5204,3400,366,5185,3302,309,5167,3185,286,5210,3083,239,5216,3066,427,5195,2919,387,5209,2812,339,5224
,5442,367,5245,5342,451,5186,5205,460,5245,5167,281,5223,5064,325,5199,4945,355,5207,4833,376,5214,4782,176,5194,4669,181,5244,4578,197,5200,4491,180,5232,4377,234,5208,4290,243,5198,4161,252,5207,4117,250,5207,3988,239,5198,3901,221,5187,3770,221,5189,3704,209,5189,3590,174,5223,3499,165,5204,3400,366,5185,3302,309,5167,3185,286,5210,3083,239,5216,3066,427,5195,2919,387,5209,2812,339,5224
,5442,367,5245,5342,451,5186,5205,460,5245,5167,281,5223,5064,325,5199,4945,355,5207,4833,376,5214,4742,400,5213,4641,376,5194,4574,396,5213,4448,405,5192,4363,432,5192,4280,439,5191,4177,450,5201,4117,427,5153,3993,422,5163,3910,396,5173,3808,418,5182,3703,403,5203,3599,407,5184,3531,376,5213,3400,366,5185,3302,309,5167,3185,286,5210,3083,239,5216,3066,427,5195,2919,387,5209,2812,339,5224
,5442,367,5245,5342,451,5186,5205,460,5245,5150,495,5213,5018,505,5192,4924,542,5172,4819,549,5182,4736,559,5210,4629,588,5181,4551,574,5200,4472,569,5228,4371,599,5163,4272,592,5163,4175,588,5163,4096,622,5200,3979,602,5163,3919,584,5172,3802,592,5172,3701,573,5209,3618,555,5181,3513,529,5172,3413,540,5182,3324,512,5182,3214,491,5182,3160,450,5184,3066,427,5195,2919,387,5209,2812,339,5224
,5391,568,5173,5323,636,5221,5195,632,5201,5121,668,5172,4997,666,5163,4887,705,5209,4788,704,5154,4723,737,5164,4629,715,5155,4535,701,5155,4513,720,5146,4358,746,5148,4264,751,5166,4171,751,5148,4096,769,5158,3984,760,5140,3909,747,5157,3795,733,5166,3719,738,5182,3621,712,5164,3525,719,5173,3422,693,5209,3354,654,5163,3240,686,5172,3165,629,5172,3074,602,5191,2974,560,5163,2836,542,5194
,5376,729,5172,5271,7409,5172,5173,765,5154,5094,825,5182,4957,817,5164,4889,857,5166,4789,878,5167,4718,865,5150,4601,896,5159,4532,866,5134,4439,875,5201,4349,874,5152,4257,906,5145,4167,913,5178,4096,902,5145,3988,889,5144,3898,885,5152,3809,883,5160,3737,890,5160,3627,888,5177,3546,846,5141,3436,856,5167,3370,815,5148,3255,816,5191,3189,793,5173,3047,789,5209,2992,747,5200,2872,704,5163
,5370,903,5173,5250,898,5191,5177,933,5175,5056,949,5150,4972,976,5159,4898,971,5160,4760,1013,5178,4687,1024,5172,4616,1016,5139,4512,1012,5155,4424,1013,5189,4334,1057,5158,4249,1041,5166,4165,1045,5175,4096,1040,5150,3993,1026,5149,3909,1050,5175,3805,1041,5134,3751,1020,5157,3594,1025,5155,3540,1017,5172,3443,979,5136,3370,979,5194,3260,980,5160,3210,940,5167,3072,926,5192,2996,879,5191,2895,880,5182
,5336,1040,5158,5210,1059,5168,5126,1084,5178,5058,1118,5172,4949,1120,5157,4870,1152,5182,4769,1136,5175,4675,1168,5162,4591,1169,5162,4494,1148,5154,4422,1187,5209,4323,1187,5149,4257,1214,5166,4161,1182,5134,4096,1189,5143,3983,1214,5152,3884,1180,5141,3816,1166,5155,3749,1150,5146,3619,1180,5178,3545,1141,5137,3453,1109,5150,3363,1104,5157,3287,1085,5148,3159,1084,5137,3095,1058,5177,2996,1045,5177,2892,1029,5184
,5319,1176,5162,5232,1203,5140,5113,1227,5182,5053,1248,5137,4942,1267,5163,4839,1265,5157,4747,1304,5152,4684,1292,5137,4587,1291,5139,4490,1297,5162,4362,1312,5141,4328,1333,5150,4252,1313,5135,4158,1319,5128,4096,1309,5135,3987,1310,5135,3893,1315,5135,3832,1318,5149,3749,1286,5139,3639,1295,5131,3562,1313,5154,3475,1290,5144,3402,1258,5180,3290,1224,5146,3180,1209,5127,3082,1184,5132,3023,1173,5172,2923,1155,5162
,5287,1295,5182,5191,1352,5178,5085,1354,5187,5041,1382,5144,4916,1409,5162,4835,1406,5149,4738,1409,5144,4684,1434,5132,4581,1414,5132,4486,1427,5127,4467,1459,5130,4317,1460,5131,4244,1445,5137,4156,1451,5131,4096,1464,5159,3962,1436,5130,3905,1468,5172,3832,1477,5159,3751,1429,5121,3648,1447,5155,3564,1408,5117,3457,1423,5159,3398,1374,5162,3281,1369,5123,3223,1342,5128,3098,1332,5178,3025,1324,5177,2903,1290,5158
,5271,1457,5128,5203,1493,5176,5054,1484,5157,5008,1523,5136,4906,1543,5163,4824,1559,5152,4748,1556,5153,4659,1551,5167,4547,1596,5153,4478,1579,5132,4404,1603,5148,4304,1620,5157,4236,1596,5111,4138,1611,5112,4081,1607,5125,3970,1593,5122,3900,1592,5148,3814,1584,5134,3742,1578,5120,3656,1585,5145,3563,1555,5162,3479,1512,5137,3406,1524,5130,3297,1474,5117,3224,1448,5135,3112,1461,5126,3031,1425,5144,2935,1405,5134
,5259,1596,5166,5207,1602,5159,5062,1596,5128,4986,1629,5153,4902,1696,5159,4817,1681,5141,4706,1717,5153,4651,1713,5146,4552,1722,5143,4458,1715,5150,4390,1711,5126,4308,1729,5135,4227,1742,5136,4149,1722,5122,4083,1721,5122,3976,1725,5122,3897,1728,5135,3831,1734,5135,3763,1724,5132,3650,1707,5117,3598,1720,5149,3489,1675,5117,3422,1644,5120,3319,1644,5123,3248,1616,5140,3118,1603,5114,3033,1556,5137,2919,1566,5149
,5233,1688,5130,5175,1743,5168,5024,1771,5155,4943,1790,5153,4888,1781,5146,4787,1830,5141,4695,1816,5136,4638,1826,5157,4540,1857,5144,4437,1848,5150,4387,1840,5109,4307,1875,5131,4220,1880,5127,4145,1902,5146,4071,1876,5127,3983,1854,5107,3909,1864,5125,3833,1862,5130,3752,1836,5114,3660,1827,5135,3601,1802,5131,3493,1799,5122,3454,1807,5135,3329,1767,5127,3256,1767,5150,3142,1744,5139,3066,1712,5162,2935,1704,5150
,5190,1844,5155,5148,1870,5132,5032,1894,5163,4961,1894,5130,4849,1931,5148,4752,1941,5140,4677,1936,5113,4627,1978,5143,4533,1950,5125,4442,1973,5128,4378,1941,5154,4294,2014,5136,4224,2026,5148,4154,2005,5136,4072,2032,5144,3989,1984,5107,3907,1987,5117,3843,1957,5102,3754,1999,5148,3660,1962,5121,3621,1948,5128,3511,1918,5112,3432,1921,5150,3338,1880,5150,3267,1877,5141,3141,1849,5122,3083,1856,5164,2961,1826,5139
,5217,1944,5149,5104,1991,5157,5009,2014,5150,4951,1966,5109,4839,2073,5150,4750,2074,5148,4665,2113,5144,4609,2100,5134,4501,2104,5143,4430,2123,5141,4362,2123,5137,4285,2112,5112,4217,2126,5114,4139,2137,5136,4074,2133,5112,3985,2114,5118,3919,2119,5118,3852,2123,5127,3770,2104,5128,3664,2092,5130,3600,2069,5116,3526,2065,5123,3444,2041,5150,3356,2007,5116,3274,1967,5130,3148,1999,5141,3086,1957,5130,2963,1949,5149
,5163,2076,5155,5066,2100,5127,5020,2112,5125,4915,2169,5146,4825,2176,5150,4739,2179,5139,4673,2205,5125,4592,2206,5117,4515,2200,5114,4422,2233,5117,4363,2272,5137,4281,2255,5122,4209,2257,5128,4148,2248,5113,4075,2274,5131,3982,2240,5117,3912,2272,5135,3850,2268,5137,3769,2227,5102,3680,2216,5126,3604,2225,5121,3516,2195,5127,3449,2133,5118,3340,2138,5120,3281,2120,5114,3183,2133,5144,3106,2087,5125,2972,2050,5114
,5149,2205,5144,5081,2204,5141,4994,2222,5122,4881,2277,5144,4811,2304,5145,4719,2305,5135,4641,2343,5143,4583,2323,5120,4487,2370,5135,4431,2352,5121,4359,2361,5123,4280,2365,5113,4208,2415,5139,4143,2402,5134,4076,2375,5116,3971,2380,5116,3920,2352,5116,3855,2378,5127,3796,2382,5143,3681,2360,5114,3624,2300,5108,3549,2337,5128,3456,2289,5132,3366,2268,5130,3285,2247,5128,3193,2211,5126,3109,2227,5144,3013,2200,5143
,5168,2314,5132,5045,2344,5148,4954,2378,5150,4869,2434,5135,4768,2412,5137,4698,2455,5137,4634,2429,5116,4560,2476,5139,4473,2475,5143,4418,2466,5134,4336,2515,5144,4264,2508,5136,4202,2511,5143,4140,2517,5148,4069,2469,5127,3987,2472,5127,3915,2488,5134,3854,2506,5139,3782,2461,5113,3691,2444,5120,3640,2437,5116,3564,2451,5140,3473,2430,5128,3361,2366,5067,3310,2380,5141,3216,2361,5123,3127,2332,5145,3014,2298,5120
,5128,2401,5118,5026,2447,5126,4933,2488,5137,4839,2522,5143,4769,2539,5141,4683,2548,5148,4620,2562,5141,4551,2572,5150,4460,2608,5140,4398,2612,5152,4323,2649,5137,4250,2649,5144,4200,2656,5141,4136,2616,5121,4071,2653,5141,3998,5553,5131,3930,2622,5127,3861,2611,5123,3779,2630,5143,3712,2600,5143,3653,2552,5131,3580,2560,5141,3493,2535,5136,3379,2531,5116,3324,2484,5123,3242,2478,5126,3132,2410,5114,3061,2419,5140
};

logic [19:0] addr;
logic [9:0] H640;
logic [8:0] V480;
logic [5:0] H36, V54;
logic [12:0] real_x, real_y, real_z;

always_comb begin
    H640 = addr % 640;
    V480 = addr / 640;
    H36 = H640 / 14;
    V54 = V480 / 12;
     
