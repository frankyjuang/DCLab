module Gaussian_Filter(
    iData,
    iStart,
    iRst,
    iClk,
    oValue,
    oDone
);

parameter bit [32:0] FIL_COEFFS [624:0] = '{
92,126,169,221,279,343,412,480,543,598,641,668,678,668,641,598,543,480,412,343,279,221,169,126,92,
126,174,233,304,384,472,566,659,747,823,882,920,933,920,882,823,747,659,566,472,384,304,233,174,126,
169,233,312,405,513,633,758,882,1000,1102,1180,1231,1247,1231,1180,1102,1000,882,758,633,513,405,312,233,169,
221,304,405,528,668,823,986,1148,1301,1433,1536,1602,1624,1602,1536,1433,1301,1148,986,823,668,528,405,304,221,
279,384,513,668,847,1042,1247,1453,1646,1814,1945,2026,2055,2026,1945,1814,1646,1453,1247,1042,847,668,513,384,279,
343,472,633,823,1042,1283,1536,1789,2026,2233,2393,2495,2530,2495,2393,2233,2026,1789,1536,1283,1042,823,633,472,343,
412,566,758,986,1247,1536,1840,2142,2427,2674,2866,2988,3029,2988,2866,2674,2427,2142,1840,1536,1247,986,758,566,412,
480,659,882,1148,1453,1789,2142,2495,2826,3115,3338,3480,3528,3480,3338,3115,2826,2495,2142,1789,1453,1148,882,659,480,
543,747,1000,1301,1646,2026,2427,2826,3202,3528,3782,3942,3997,3942,3782,3528,3202,2826,2427,2026,1646,1301,1000,747,543,
598,823,1102,1433,1814,2233,2674,3115,3528,3888,4167,4344,4404,4344,4167,3888,3528,3115,2674,2233,1814,1433,1102,823,598,
641,882,1180,1536,1945,2393,2866,3338,3782,4167,4465,4655,4720,4655,4465,4167,3782,3338,2866,2393,1945,1536,1180,882,641,
668,920,1231,1602,2026,2495,2988,3480,3942,4344,4655,4852,4920,4852,4655,4344,3942,3480,2988,2495,2026,1602,1231,920,668,
678,933,1247,1624,2055,2530,3029,3528,3997,4404,4720,4920,4989,4920,4720,4404,3997,3528,3029,2530,2055,1624,1247,933,678,
668,920,1231,1602,2026,2495,2988,3480,3942,4344,4655,4852,4920,4852,4655,4344,3942,3480,2988,2495,2026,1602,1231,920,668,
641,882,1180,1536,1945,2393,2866,3338,3782,4167,4465,4655,4720,4655,4465,4167,3782,3338,2866,2393,1945,1536,1180,882,641,
598,823,1102,1433,1814,2233,2674,3115,3528,3888,4167,4344,4404,4344,4167,3888,3528,3115,2674,2233,1814,1433,1102,823,598,
543,747,1000,1301,1646,2026,2427,2826,3202,3528,3782,3942,3997,3942,3782,3528,3202,2826,2427,2026,1646,1301,1000,747,543,
480,659,882,1148,1453,1789,2142,2495,2826,3115,3338,3480,3528,3480,3338,3115,2826,2495,2142,1789,1453,1148,882,659,480,
412,566,758,986,1247,1536,1840,2142,2427,2674,2866,2988,3029,2988,2866,2674,2427,2142,1840,1536,1247,986,758,566,412,
343,472,633,823,1042,1283,1536,1789,2026,2233,2393,2495,2530,2495,2393,2233,2026,1789,1536,1283,1042,823,633,472,343,
279,384,513,668,847,1042,1247,1453,1646,1814,1945,2026,2055,2026,1945,1814,1646,1453,1247,1042,847,668,513,384,279,
221,304,405,528,668,823,986,1148,1301,1433,1536,1602,1624,1602,1536,1433,1301,1148,986,823,668,528,405,304,221,
169,233,312,405,513,633,758,882,1000,1102,1180,1231,1247,1231,1180,1102,1000,882,758,633,513,405,312,233,169,
126,174,233,304,384,472,566,659,747,823,882,920,933,920,882,823,747,659,566,472,384,304,233,174,126,
92,126,169,221,279,343,412,480,543,598,641,668,678,668,641,598,543,480,412,343,279,221,169,126,92
};
parameter IDLE  =   1'b0;
parameter CALC  =   1'b1;

input       [9:0]   iData   [624:0];
input               iStart;
input               iRst;
input               iClk;
output reg          oValue;
output reg          oDone;

logic   [1:0]   state_r, state_w;
logic   [9:0]   counter_r, counter_w;
logic   [39:0]  sum_r, sum_w;
logic   [9:0]   value_r, value_w;
logic           done_r, done_w;

assign oValue   =   value_r;
assign oDone    =   done_r;

always_comb begin
    state_w = state_r;
    counter_w = counter_r;
    sum_w = sum_r;
    value_w = value_r;
    done_w = done_r;
    case(state_r)
        IDLE:
            begin
                done_w = 0;
                if (iStart) begin
                    state_w = CALC;
                    counter_w = 0;
                    sum_w = 0;
                end
            end
        CALC:
            begin
                for (counter_w=1; counter_w < 625; counter_w=counter_w+1) begin
                    sum_w = sum_w + FIL_COEFFS[counter_w] * iData[counter_w];
                end
                state_w = IDLE;
                done_w = 1;
                value_w = (sum_w >> 20);
                /*
                if (counter_r < 625) begin
                    sum_w = sum_r + FIL_COEFFS[counter_r] * iData[counter_r];
                    counter_r = counter_w + 1;
                end
                if (counter_r == 624) begin
                    state_w = IDLE;
                    done_w = 1;
                    value_w = (sum_r >> 20);
                end
                */
            end
    endcase
end

always_ff@(posedge iClk or negedge iRst) begin
    if(!iRst) begin
        state_r     <=  IDLE;
        counter_r   <=  0;
        sum_r       <=  0;
        value_r     <=  0;
        done_r      <=  0;
    end else begin
        state_r     <=  state_w;
        counter_r   <=  counter_w;
        sum_r       <=  sum_w;
        value_r     <=  value_w;
        done_r      <=  done_w;
    end
end

endmodule
